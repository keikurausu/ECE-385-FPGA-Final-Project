//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Viral Mehta                                                        --
//    Spring 2005                                                        --
//                                                                       --
//    Modified by Stephen Kempf 03-01-2006                               --
//                              03-12-2007                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 298 Lab 7                                         --
//    UIUC ECE Department                                                --
//-------------------------------------------------------------------------


module  ball2 ( input Reset, frame_clk, press,
					input [7:0] keycode,
               output [9:0]  BallX, BallY, BallS );
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion, Ball_Size;
	 
    parameter [9:0] Ball_X_Center=160;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center=240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min=0;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max=639;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min=0;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max=479;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step=1;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step=1;      // Step size on the Y axis

    assign Ball_Size = 4;  // assigns the value 4 as a 10-digit binary number, ie "0000000100"
   
    always_ff @ (posedge Reset or posedge frame_clk )
    begin: Move_Ball
        if (Reset)  // Asynchronous Reset
        begin 
            Ball_Y_Motion <= 10'd0; //Ball_Y_Step;
				Ball_X_Motion <= 10'd0; //Ball_X_Step;
				Ball_Y_Pos <= Ball_Y_Center;
				Ball_X_Pos <= Ball_X_Center;
        end
           
        else 
		  
		  begin 
		  if ( (Ball_Y_Pos + Ball_Size) >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
					  Ball_Y_Motion <= (~ (Ball_Y_Step) + 1'b1);  // 2's complement.
					  
				 else if ( (Ball_Y_Pos - Ball_Size) <= Ball_Y_Min )  // Ball is at the top edge, BOUNCE!
					  Ball_Y_Motion <= Ball_Y_Step;
					
				 else 
					  Ball_Y_Motion <= Ball_Y_Motion;  // Ball is somewhere in the middle, don't bounce, just keep moving
					 
				
				if ( (Ball_X_Pos + Ball_Size) >= Ball_X_Max)
					 Ball_X_Motion <= (~ (Ball_X_Step) + 1'b1);
					
					
				else if ( (Ball_X_Pos - Ball_Size) <= Ball_X_Min)
					 Ball_X_Motion <=Ball_X_Step;
				else
					Ball_X_Motion <= Ball_X_Motion;
					
				
			
			case(keycode)
			8'h43: //W ps/2
				begin
				if(press == 1'b1)
					begin
					Ball_Y_Motion <= -1;
					Ball_X_Motion <= 0;
					end
				end
			8'h3B: //A ps/2
				begin
					if(press == 1'b1)
					begin
					Ball_Y_Motion <= 0;
					Ball_X_Motion <= -1;
					end
				end
			8'h42: //S ps/2
				begin
					if(press == 1'b1)
					begin
					Ball_X_Motion <= 0;
					Ball_Y_Motion <= 1;
					end
				end
			8'h4B: //D ps/2
				begin
					if(press == 1'b1)
					begin
					Ball_X_Motion <= 1;
					Ball_Y_Motion <= 0;
					end
				end
			default: ;
			 endcase
			begin
			
			if ( (Ball_Y_Pos + Ball_Size) >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
			begin
					  Ball_Y_Motion <= (~ (Ball_Y_Step) + 1'b1);  // 2's complement.
					  
					  end
				 else if ( (Ball_Y_Pos - Ball_Size) <= Ball_Y_Min )  // Ball is at the top edge, BOUNCE!
				 begin
					  Ball_Y_Motion <= Ball_Y_Step;
					  
					  end
				 
				 
				// Ball_X_Motion <= Ball_X_Motion;  // You need to remove this and make both X and Y respond to keyboard input
				
				if ( (Ball_X_Pos + Ball_Size) >= Ball_X_Max)
				begin
					 Ball_X_Motion <= (~ (Ball_X_Step) + 1'b1);
					
					 end
				else if ( (Ball_X_Pos - Ball_Size) <= Ball_X_Min)
				begin
					 Ball_X_Motion <=Ball_X_Step;
					 
				end

				
			end
			
		 
		  
				  Ball_Y_Pos <= (Ball_Y_Pos + Ball_Y_Motion);  // Update ball position
				 Ball_X_Pos <= (Ball_X_Pos + Ball_X_Motion);
			
				
	  
		end
		
    end
       
    assign BallX = Ball_X_Pos;
   
    assign BallY = Ball_Y_Pos;
   
    assign BallS = Ball_Size;
    

endmodule
